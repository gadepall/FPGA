module sevenseg(output reg a, output reg b, output reg c, output reg d,output reg e, output reg f,output reg g);
    initial
    begin
    a=0;
    b=0;
    c=0;
    d=0;
    e=0;
    f=0;
    g=1;
    end
endmodule
