//Program for turning LED on and off
module example(output reg A);

//  reg[26:0] delay;
//wire A;
//  always@(posedge clk) 
	initial
	begin
//  delay = delay+1;
//  if(delay==27'b101111101011110000100000000) begin
 //  delay =27'b0;
	A=1;
	end
//   end
endmodule
