module display_decoder(

input wire A,
input wire B,
input wire C,
input wire D,

output reg a,
output reg b,
output reg c,
output reg d);



assign a=A;
assign b=B;
assign c=C;
assign d=D;
endmodule
