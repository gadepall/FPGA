`timescale 1ns / 1ps
///////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 31.10.2017 14:17:14
// Design Name: 
// Module Name: sevenseg
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
/////////////////////


module sevenseg(input wire clk, output reg a, output reg b, output reg c, output reg d,output reg e, output reg f,output reg g 

    );
    initial
    begin
    a=1;
    b=0;
    c=0;
    d=1;
    e=1;
    f=1;
    g=1;
    end
endmodule
